-- $Id: $
-- File name:   rkeyGen.vhd
-- Created:     4/10/2011
-- Author:      Samuel Oshin
-- Lab Section: 337-02
-- Version:     1.0  Initial Design Entry
-- Description: ROUND KEY GENERATORRRRRRR!!!@!@!@!@!


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

