-- $Id: $
-- File name:   B_SRAM1.vhd
-- Created:     4/10/2011
-- Author:      Yonatan Feleke
-- Lab Section: 337-02
-- Version:     1.0  Initial Design Entry
-- Description: this is a wrapper that will contain an sram. Will strore prvalues.


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

