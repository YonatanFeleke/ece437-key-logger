-- $Id: $
-- File name:   edge_detect.vhd
-- Created:     2/21/2011
-- Author:      Brian Crone
-- Lab Section: 337-02
-- Version:     1.0  Initial Design Entry
-- Description: Source code for Edge_detect for the USB receiver.


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

Entity U_EDGE_DETECT is
	port(D_CLK	:	in	std_logic;
			 rst_n	:	in	std_logic;
			 d_plus	:	in	std_logic;
			 d_edge	:	out	std_logic);
	end U_EDGE_DETECT;

architecture behavioral of U_EDGE_DETECT is
	signal current, previous : std_logic;
	begin
		detect	:	process(D_CLK, rst_n)
		begin
			--current <= D_PLUS;
			if(rst_n = '1') then
				D_EDGE <= '0';
				current <= '1';
				previous <= '1';
			elsif(rising_edge(D_CLK)) then
				current <= D_PLUS;
				previous <= current;
				if (current = '1' and previous = '0') or (current = '0' and previous = '1') then
					D_EDGE <= '1';
				else D_EDGE <= '0';
				end if;
			end if;
		end process detect;
	
end behavioral;
			

