-- $Id: $
-- File name:   B_RCU.vhd
-- Created:     4/10/2011
-- Author:      Yonatan Feleke
-- Lab Section: 337-02
-- Version:     1.0  Initial Design Entry
-- Description: Control unit for sram and enabling bluetoot coding


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

