-- $Id: $
-- File name:   B_Header.vhd
-- Created:     4/10/2011
-- Author:      Yonatan Feleke
-- Lab Section: 337-02
-- Version:     1.0  Initial Design Entry
-- Description: Outputs the header on the bus to sram


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

